package data_types_pkg is
	type username_array_of_8_characters is array (1 to 8) of character;
	type password_array_of_4_characters is array (1 to 4) of character;
end package data_types_pkg;